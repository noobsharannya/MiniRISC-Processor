module comp_less(input[31:0] a,output res);
    assign res=input[31];
endmodule